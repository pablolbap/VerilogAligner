include "machin"
include   "machin2"
include     "machin3

wire [6:0]   truc     = 0;
;

wire   [25:0] mac   = 1;


assign truc2 = truc[0];
